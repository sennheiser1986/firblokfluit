Package Constants_pack is

	constant Threshold       : real    := 0.0001;
	constant SampleFrequency : integer := 44100;
	constant ClockFrequency  : integer := 100000000;
	
end Constants_pack;

package body Constants_pack is
end Constants_pack;