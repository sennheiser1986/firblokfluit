library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


Package Constants_pack is

	constant Threshold       : integer := 3;
	constant SampleFrequency : integer := 48000;
	constant ClockFrequency  : integer := 100000000;
	
end Constants_pack;

package body Constants_pack is
end Constants_pack;